library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity amp_lock is
		Port ( clk 		: in  STD_LOGIC;
			   reset 	: in  STD_LOGIC;
			   comp_state : in STD_LOGIC;
			   saw_amp 	: in integer;
			   locked_amp: out std_logic_vector (10 downto 0)
			 );
end amp_lock;

architecture Behavioral of amp_lock is

signal  i_comp_state: std_logic;
signal  lastState: std_logic;
signal  i_locked_amp: integer;--std_logic_vector (10 downto 0);
--signal  table_output : std_logic_vector (8 downto 0);

type test is array (0 to 2047) of integer;--std_logic_vector(8 downto 0);
--signal distance: test := ("100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100100111", "100100111", "100100010", "100011101", "100011000", "100010011", "100001110", "100001110", "100001110", "100001001", "100000100", "100000100", "011111111", "011111010", "011110101", "011110000", "011110000", "011101011", "011101011", "011100110", "011100110", "011100001", "011100001", "011011100", "011011100", "011010111", "011010111", "011010010", "011010010", "011010010", "011001101", "011001101", "011001101", "011001000", "011001000", "011001000", "011000011", "011000011", "011000011", "011000011", "010111110", "010111110", "010111110", "010111001", "010111001", "010111001", "010110100", "010110100", "010110100", "010101111", "010101111", "010101111", "010101010", "010101010", "010101010", "010100101", "010100101", "010100101", "010100000", "010100000", "010100000", "010011011", "010011011", "010011011", "010011011", "010011011", "010011011", "010010110", "010010110", "010010110", "010010001", "010010001", "010010001", "010001100", "010001100", "010001100", "010001100", "010001100", "010001100", "010000111", "010000111", "010000111", "010000010", "010000010", "010000010", "001111101", "001111101", "001111101", "001111101", "001111101", "001111101", "001111000", "001111000", "001111000", "001111000", "001111000", "001111000", "001110011", "001110011", "001110011", "001110011", "001110011", "001110011", "001101110", "001101110", "001101110", "001101110", "001101110", "001101110", "001101001", "001101001", "001101001", "001101001", "001101001", "001101001", "001101001", "001101001", "001100100", "001100100", "001100100", "001100100", "001100100", "001100100", "001100100", "001100100", "001100100", "001011111", "001011111", "001011111", "001011111", "001011111", "001011111", "001011111", "001011111", "001011111", "001011010", "001011010", "001011010", "001011010", "001011010", "001011010", "001011010", "001011010", "001011010", "001011010", "001011010", "001011010", "001010101", "001010101", "001010101", "001010101", "001010101", "001010101", "001010101", "001010101", "001010101", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110");
signal distance: test := (300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 290, 280, 280, 280, 280, 280, 280, 280, 280, 280, 280, 280, 280, 270, 270, 270, 270, 270, 270, 270, 270, 270, 270, 270, 270, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 260, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 250, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 220, 220, 220, 220, 220, 220, 220, 220, 220, 220, 220, 220, 210, 210, 210, 210, 210, 210, 210, 210, 210, 210, 210, 210, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 190, 190, 190, 190, 190, 190, 190, 190, 190, 190, 190, 190, 190, 190, 190, 190, 190, 190, 180, 180, 180, 180, 180, 180, 180, 180, 180, 180, 180, 180, 180, 180, 180, 180, 180, 180, 175, 175, 175, 175, 175, 175, 175, 175, 175, 175, 175, 175, 175, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 165, 165, 165, 165, 165, 165, 165, 165, 165, 165, 165, 165, 160, 160, 160, 160, 160, 160, 160, 160, 160, 160, 160, 160, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 150, 150, 150, 150, 150, 150, 150, 150, 150, 150, 150, 150, 150, 150, 150, 150, 150, 150, 145, 145, 145, 145, 145, 145, 145, 145, 145, 145, 145, 145, 145, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30);
	
begin

process(clk, reset, i_comp_state)
begin
	if (reset = '1') then					
        i_locked_amp <= 0;--"00000000000";
        lastState <= i_comp_state;
        
    elsif(rising_edge(clk)) then
        if(lastState = '1' and i_comp_state = '0') then      
             i_locked_amp <= saw_amp;--std_logic_vector(to_unsigned(saw_amp, 11));
	    end if;
        lastState <= i_comp_state;
    end if;
end process;

locked_amp <= std_logic_vector(to_unsigned(distance(i_locked_amp), 11));--i_locked_amp;
i_comp_state <= comp_state;

end Behavioral;
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity amp_lock is
		Port ( clk 		: in  STD_LOGIC;
			   reset 	: in  STD_LOGIC;
			   comp_state : in STD_LOGIC;
			   saw_amp 	: in integer;
			   locked_amp: out std_logic_vector (8 downto 0)
			 );
end amp_lock;

architecture Behavioral of amp_lock is

signal  i_comp_state: std_logic;
signal  lastState: std_logic;
signal  i_locked_amp: integer;--std_logic_vector (8 downto 0);
--signal  table_output : std_logic_vector (8 downto 0);

type test is array (511 downto 0) of integer;--std_logic_vector(8 downto 0);
--signal distance: test := ("100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100101100", "100100111", "100100111", "100100010", "100011101", "100011000", "100010011", "100001110", "100001110", "100001110", "100001001", "100000100", "100000100", "011111111", "011111010", "011110101", "011110000", "011110000", "011101011", "011101011", "011100110", "011100110", "011100001", "011100001", "011011100", "011011100", "011010111", "011010111", "011010010", "011010010", "011010010", "011001101", "011001101", "011001101", "011001000", "011001000", "011001000", "011000011", "011000011", "011000011", "011000011", "010111110", "010111110", "010111110", "010111001", "010111001", "010111001", "010110100", "010110100", "010110100", "010101111", "010101111", "010101111", "010101010", "010101010", "010101010", "010100101", "010100101", "010100101", "010100000", "010100000", "010100000", "010011011", "010011011", "010011011", "010011011", "010011011", "010011011", "010010110", "010010110", "010010110", "010010001", "010010001", "010010001", "010001100", "010001100", "010001100", "010001100", "010001100", "010001100", "010000111", "010000111", "010000111", "010000010", "010000010", "010000010", "001111101", "001111101", "001111101", "001111101", "001111101", "001111101", "001111000", "001111000", "001111000", "001111000", "001111000", "001111000", "001110011", "001110011", "001110011", "001110011", "001110011", "001110011", "001101110", "001101110", "001101110", "001101110", "001101110", "001101110", "001101001", "001101001", "001101001", "001101001", "001101001", "001101001", "001101001", "001101001", "001100100", "001100100", "001100100", "001100100", "001100100", "001100100", "001100100", "001100100", "001100100", "001011111", "001011111", "001011111", "001011111", "001011111", "001011111", "001011111", "001011111", "001011111", "001011010", "001011010", "001011010", "001011010", "001011010", "001011010", "001011010", "001011010", "001011010", "001011010", "001011010", "001011010", "001010101", "001010101", "001010101", "001010101", "001010101", "001010101", "001010101", "001010101", "001010101", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001010000", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001001011", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000110", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "001000001", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000111100", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110111", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000110010", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101101", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000101000", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000100011", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110", "000011110");
signal distance: test := (30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 85, 85, 85, 85, 85, 85, 85, 85, 85, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 95, 95, 95, 95, 95, 95, 95, 95, 95, 100, 100, 100, 100, 100, 100, 100, 100, 100, 105, 105, 105, 105, 105, 105, 105, 105, 110, 110, 110, 110, 110, 110, 115, 115, 115, 115, 115, 115, 120, 120, 120, 120, 120, 120, 125, 125, 125, 125, 125, 125, 130, 130, 130, 135, 135, 135, 140, 140, 140, 140, 140, 140, 145, 145, 145, 150, 150, 150, 155, 155, 155, 155, 155, 155, 160, 160, 160, 165, 165, 165, 170, 170, 170, 175, 175, 175, 180, 180, 180, 185, 185, 185, 190, 190, 190, 195, 195, 195, 195, 200, 200, 200, 205, 205, 205, 210, 210, 210, 215, 215, 220, 220, 225, 225, 230, 230, 235, 235, 240, 240, 245, 250, 255, 260, 260, 265, 270, 270, 270, 275, 280, 285, 290, 295, 295, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300, 300);
	
begin

process(clk, reset, i_comp_state)
begin
	if (reset = '1') then					
        i_locked_amp <= 0;--"000000000";
        lastState <= i_comp_state;
        
    elsif(rising_edge(clk)) then
        if(lastState = '1' and i_comp_state = '0') then      
             i_locked_amp <= saw_amp;--std_logic_vector(to_unsigned(saw_amp, 9));
	    end if;
        lastState <= i_comp_state;
    end if;
end process;

locked_amp <= std_logic_vector(to_unsigned(distance(i_locked_amp), 9));
i_comp_state <= comp_state;

end Behavioral;